*Inverter simulation

.lib "~/software/PDKs/sky130A/libs.tech/ngspice/sky130.lib.spice" tt

Xinv Y A VPWR VGND VGND VPWR inverter

.subckt inverter Y A NWELL VSUBS VGND VPWR
X0 Y A VPWR NWELL sky130_fd_pr__pfet_01v8 ad=6e+11p pd=3.2e+06u as=5.5e+11p ps=3.1e+06u w=1e+06u l=150000u
X1 Y A VGND VSUBS sky130_fd_pr__nfet_01v8 ad=6e+11p pd=3.2e+06u as=5.5e+11p ps=3.1e+06u w=650000u l=150000u
.ends

*set gnd and power
Vgnd VGND 0 0
Vdd VPWR VGND 1.8

*create pulse
Vin A VGND pulse(0 1.8 1p 10p 10p 1n 3n)
.tran 10e-12 2e-09 0e-00

.control
run
set color0 = white
set color1 = black
plot A Y
plot VPWR
.endc

.end


