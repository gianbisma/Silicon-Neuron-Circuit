magic
tech sky130A
timestamp 1686368637
<< nwell >>
rect -130 145 320 285
<< nmos >>
rect 0 -40 15 60
rect 225 -40 240 60
rect 0 -231 15 -131
rect 225 -231 240 -131
<< pmos >>
rect 0 165 15 265
rect 225 165 240 265
<< ndiff >>
rect -55 45 0 60
rect -55 -25 -40 45
rect -15 -25 0 45
rect -55 -40 0 -25
rect 15 45 75 60
rect 15 -25 30 45
rect 55 -25 75 45
rect 15 -40 75 -25
rect 170 45 225 60
rect 170 -25 185 45
rect 210 -25 225 45
rect 170 -40 225 -25
rect 240 45 300 60
rect 240 -25 255 45
rect 280 -25 300 45
rect 240 -40 300 -25
rect -55 -146 0 -131
rect -55 -216 -40 -146
rect -15 -216 0 -146
rect -55 -231 0 -216
rect 15 -146 75 -131
rect 15 -216 30 -146
rect 55 -216 75 -146
rect 15 -231 75 -216
rect 170 -146 225 -131
rect 170 -216 185 -146
rect 210 -216 225 -146
rect 170 -231 225 -216
rect 240 -146 300 -131
rect 240 -216 255 -146
rect 280 -216 300 -146
rect 240 -231 300 -216
<< pdiff >>
rect -55 250 0 265
rect -55 180 -40 250
rect -15 180 0 250
rect -55 165 0 180
rect 15 250 75 265
rect 15 180 30 250
rect 55 180 75 250
rect 15 165 75 180
rect 170 250 225 265
rect 170 180 185 250
rect 210 180 225 250
rect 170 165 225 180
rect 240 250 300 265
rect 240 180 255 250
rect 280 180 300 250
rect 240 165 300 180
<< ndiffc >>
rect -40 -25 -15 45
rect 30 -25 55 45
rect 185 -25 210 45
rect 255 -25 280 45
rect -40 -216 -15 -146
rect 30 -216 55 -146
rect 185 -216 210 -146
rect 255 -216 280 -146
<< pdiffc >>
rect -40 180 -15 250
rect 30 180 55 250
rect 185 180 210 250
rect 255 180 280 250
<< psubdiff >>
rect -110 45 -55 60
rect -110 -25 -95 45
rect -70 -25 -55 45
rect -110 -40 -55 -25
rect 115 45 170 60
rect 115 -25 130 45
rect 155 -25 170 45
rect 115 -40 170 -25
rect -110 -146 -55 -131
rect -110 -216 -95 -146
rect -70 -216 -55 -146
rect -110 -231 -55 -216
rect 115 -146 170 -131
rect 115 -216 130 -146
rect 155 -216 170 -146
rect 115 -231 170 -216
<< nsubdiff >>
rect -110 250 -55 265
rect -110 180 -95 250
rect -70 180 -55 250
rect -110 165 -55 180
rect 115 250 170 265
rect 115 180 130 250
rect 155 180 170 250
rect 115 165 170 180
<< psubdiffcont >>
rect -95 -25 -70 45
rect 130 -25 155 45
rect -95 -216 -70 -146
rect 130 -216 155 -146
<< nsubdiffcont >>
rect -95 180 -70 250
rect 130 180 155 250
<< poly >>
rect 45 310 85 320
rect 45 295 55 310
rect 0 290 55 295
rect 75 295 85 310
rect 75 290 240 295
rect 0 280 240 290
rect 0 265 15 280
rect 225 265 240 280
rect 0 150 15 165
rect 225 150 240 165
rect -25 105 15 115
rect -25 85 -15 105
rect 5 85 15 105
rect -25 75 15 85
rect 200 105 240 115
rect 200 85 210 105
rect 230 85 240 105
rect 200 75 240 85
rect 0 60 15 75
rect 225 60 240 75
rect 0 -55 15 -40
rect 225 -55 240 -40
rect 45 -90 85 -80
rect 45 -100 55 -90
rect 0 -110 55 -100
rect 75 -110 85 -90
rect 0 -120 85 -110
rect 0 -131 15 -120
rect 225 -131 240 -115
rect 0 -246 15 -231
rect 225 -246 240 -231
<< polycont >>
rect 55 290 75 310
rect -15 85 5 105
rect 210 85 230 105
rect 55 -110 75 -90
<< locali >>
rect 45 310 85 320
rect 45 290 55 310
rect 75 290 85 310
rect 45 280 85 290
rect 45 260 65 280
rect -105 250 -5 260
rect -105 180 -95 250
rect -70 180 -40 250
rect -15 180 -5 250
rect -105 170 -5 180
rect 20 250 65 260
rect 20 180 30 250
rect 55 180 65 250
rect 20 170 65 180
rect 120 250 220 260
rect 120 180 130 250
rect 155 180 185 250
rect 210 180 220 250
rect 120 170 220 180
rect 245 250 290 260
rect 245 180 255 250
rect 280 180 290 250
rect 245 170 290 180
rect -130 105 15 115
rect -130 95 -15 105
rect -25 85 -15 95
rect 5 85 15 105
rect -25 75 15 85
rect 45 55 65 170
rect 95 105 240 115
rect 95 95 210 105
rect 200 85 210 95
rect 230 85 240 105
rect 200 75 240 85
rect 270 55 290 170
rect -105 45 -5 55
rect -105 -25 -95 45
rect -70 -25 -40 45
rect -15 -25 -5 45
rect -105 -35 -5 -25
rect 20 45 65 55
rect 20 -25 30 45
rect 55 -25 65 45
rect 20 -35 65 -25
rect 120 45 220 55
rect 120 -25 130 45
rect 155 -25 185 45
rect 210 -25 220 45
rect 120 -35 220 -25
rect 245 45 290 55
rect 245 -25 255 45
rect 280 -25 290 45
rect 245 -35 290 -25
rect 45 -80 65 -35
rect 45 -90 85 -80
rect 45 -110 55 -90
rect 75 -110 85 -90
rect 45 -120 85 -110
rect 45 -136 65 -120
rect 270 -136 290 -35
rect -105 -146 -5 -136
rect -105 -216 -95 -146
rect -70 -216 -40 -146
rect -15 -216 -5 -146
rect -105 -226 -5 -216
rect 20 -146 65 -136
rect 20 -216 30 -146
rect 55 -216 65 -146
rect 20 -226 65 -216
rect 120 -146 220 -136
rect 120 -216 130 -146
rect 155 -216 185 -146
rect 210 -216 220 -146
rect 120 -226 220 -216
rect 245 -146 290 -136
rect 245 -216 255 -146
rect 280 -216 290 -146
rect 245 -226 290 -216
<< viali >>
rect -95 180 -70 250
rect -40 180 -15 250
rect 130 180 155 250
rect 185 180 210 250
rect -95 -25 -70 45
rect -40 -25 -15 45
rect 130 -25 155 45
rect 185 -25 210 45
rect -95 -216 -70 -146
rect -40 -216 -15 -146
rect 130 -216 155 -146
rect 185 -216 210 -146
<< metal1 >>
rect -130 250 320 260
rect -130 180 -95 250
rect -70 180 -40 250
rect -15 180 130 250
rect 155 180 185 250
rect 210 180 320 250
rect -130 170 320 180
rect 45 165 70 170
rect -130 45 320 55
rect -130 -25 -95 45
rect -70 -25 -40 45
rect -15 -25 130 45
rect 155 -25 185 45
rect 210 -25 320 45
rect -130 -35 320 -25
rect -130 -146 320 -136
rect -130 -216 -95 -146
rect -70 -216 -40 -146
rect -15 -216 130 -146
rect 155 -216 185 -146
rect 210 -216 320 -146
rect -130 -226 320 -216
<< labels >>
rlabel metal1 -130 170 -95 260 1 VPWR
port 5 n
rlabel metal1 -130 -226 -95 -136 1 VGND
port 6 n
rlabel polycont -15 85 5 105 1 V
port 3 n
rlabel polycont 210 85 230 105 1 Vth
port 4 n
rlabel locali 45 45 65 180 1 VB
port 1 n
rlabel locali 270 45 290 180 1 VA
port 2 n
rlabel poly 225 -131 240 -115 1 Vbias
port 7 n
<< end >>
